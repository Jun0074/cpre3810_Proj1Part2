library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IFID_Register is
  generic (
    N : integer := 32  -- width of PC and instruction
  );
  port (
    i_CLK     : in  std_logic;
    i_RST     : in  std_logic;                 -- synchronous reset (active high)
    i_FLUSH   : in  std_logic;                 -- insert bubble/NOP this cycle (active high)

    -- inputs from IF stage
    i_PC      : in  std_logic_vector(N-1 downto 0);
    i_Instr   : in  std_logic_vector(31 downto 0);

    -- outputs to ID stage
    o_PC      : out std_logic_vector(N-1 downto 0);
    o_Instr   : out std_logic_vector(31 downto 0)
  );
end IFID_Register;

architecture structure of IFID_Register is

  -- For RISC-V, NOP = ADDI x0, x0, 0 = 0x00000013
  constant NOP_32 : std_logic_vector(31 downto 0) := x"00000013";

  signal s_holding_PC : std_logic_vector(N-1 downto 0);
  signal s_holding_Instr        : std_logic_vector(31 downto 0);

begin
  process(iCLK)
  begin
    if rising_edge(iCLK) then
      if iRST = '1' then
	-- Reset holding values
        s_holding_PC      <= (others => '0'); -- Set PC to 0 until no longer reset
        s_holding_Instr   <= NOP_32;

      elsif iFLUSH = '1' then
        -- Convert the next ID stage cycle into a bubble (Don't update holding PC value)
        s_holding_Instr   <= NOP_32;
      
      else
        -- Normal pipeline advance
        s_holding_PC      <= i_PC;
        s_holding_Instr   <= i_Instr;

      end if;
    end if;
  end process;

  -- Update output with holding signals
  o_PC      <= s_holding_PC;
  o_Instr   <= s_holding_Instr;

end structure;
